19D070052 Sheel Shah Solar IV
.include Solar_Cell.txt

r1 0 21 100
x1 21 31 solar_cell IL_val = 8e-3 rsh_val = 100
v_dummy1 0 31 0

r2 0 22 100
x2 22 32 solar_cell IL_val = 8e-3 rsh_val = 500
v_dummy2 0 32 0

r3 0 23 100
x3 23 33 solar_cell IL_val = 8e-3 rsh_val = 5k
v_dummy3 0 33 0

* start control
.control
set color0 = rgb:f/f/e
set color1 = rgb:1/1/1

run

dc r1 1 500 1
let i1 = i(v_dummy1)
let v1 = v(21)-v(31)
let p1 = i1*v1

dc r2 1 500 1
let i2 = i(v_dummy2)
let v2 = v(22)-v(32)
let p2 = i2*v2

dc r3 1 500 1
let i3 = i(v_dummy3)
let v3 = v(23)-v(33)
let p3 = i3*v3

plot dc1.i1 vs dc1.v1, dc2.i2 vs dc2.v2, dc3.i3 vs dc3.v3
plot dc1.p1 vs dc1.v1, dc2.p2 vs dc2.v2, dc3.p3 vs dc3.v3

** values(rs 0 10 30)
** i_sc = 8m, 7.9m, 7.6m
** v_oc = 0.42, 0.41, 0.39
** p_mp = 2.16m, 1.74m, 1.12m
** ff = 0.64, 0.54, 0.38

** values(rsh 100 500 5k)
** i_sc = 7.2m, 7.8m, 8m
** v_oc = 0.38, 0.41, 0.42
** p_mp = 1.11m, 1.66m, 1.80m
** ff = 0.41, 0.52, 0.54

* end control
.endc

.end