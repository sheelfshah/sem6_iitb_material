Sheel Shah 19D070052

.include bc547.txt

q0 0 1 2 bc547a
r2 3 2 100
i_source 0 1
v_ce 3 0 

.dc v_ce 0 100 0.1 i_source 0 1m 0.1m
.control
run

plot -i(v_ce) vs v(2)

.endc
.end 
