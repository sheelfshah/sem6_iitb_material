19D070052 Sheel Shah I_d vs V_ds

.include ALD1105N.txt

** 1 2 3 4: drain gate source body
m1 1 2 0 4 ALD1105N
v_dd 4 0 0
v_id 10 1 0
v_ds 10 0 5
v_gs 2 0


.dc v_gs 0 5 0.1

* start control
.control
set color0 = rgb:f/f/e
set color1 = rgb:1/1/1

run

plot (i(v_id)) vs v(2)

** v_t by linear region's intercept: 0.706
** K = 2 * slope * slope = 5.107080e-04 A/V^2
.endc

.end