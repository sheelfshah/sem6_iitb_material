19D070052 Sheel Shah Solar IV
.include Solar_Cell.txt

v_dc 1 0

r1 1 21 100
x1 21 31 solar_cell IL_val = 0e-3
v_dummy1 31 0 0

r2 1 22 100
x2 22 32 solar_cell IL_val = 8e-3
v_dummy2 32 0 0

r3 1 23 100
x3 23 33 solar_cell IL_val = 10e-3
v_dummy3 33 0 0
** 1: dark, 2: 8mA, 3: 10mA
.dc v_dc 0.5 2 0.01

* start control
.control
set color0 = rgb:f/f/e
set color1 = rgb:1/1/1

run

plot log(i(v_dummy1)) vs v(21)-v(31), log(i(v_dummy2)) vs v(22)-v(32), log(i(v_dummy3)) vs v(23)-v(33)
* plot i(v_dummy1) vs v(21)-v(31), i(v_dummy2) vs v(22)-v(32), i(v_dummy3) vs v(23)-v(33)
** dx/dy: 0.152159, 0.136435, 0.121013
** eta = (dx/dy)/V_t = 3.89, 3.27, 2.69


* end control
.endc

.end