19D070052 Sheel Shah I_d vs V_ds

.include PMOS_NMOS.txt

** 1 2 0 4: drain gate source body
m1 1 2 5 4 cmosp L=0.4u W=4u
v_dd 4 0 3.3
v_id 10 1 0
v_ds 10 0
v_gs 2 0 -3.3
r_l 5 0 10k


.dc v_ds -3.3 3.3 0.01

* start control
.control
set color0 = rgb:f/f/e
set color1 = rgb:1/1/1

run

plot v(5) vs v(10)
plot abs(v(10)/i(v_id))-10k vs v(10)


.endc

.end

** pmos has hgher r due to higher v_th
