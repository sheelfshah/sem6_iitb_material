19D070052 Sheel Shah I_d vs V_ds

.include NMOSFET.txt

** 1 2 3 4: drain gate source body
m1 1 2 0 4 NMOSFET W=30u L=0.4u
v_dd 4 0 0
v_id 10 1 0
v_ds 10 0 0.3
v_gs 2 0


.dc v_gs 0 3.3 0.01 temp 25 125 50

* start control
.control
run
 
plot log10(i(v_id)) vs v(2)

** ss: 25: 98.7, 75: 111.6, 125: 126.0 (mV/dec)
** off current: 6.3e-12, 6.3e-11, 3.2e-10

.endc

.end