19D070052 Sheel Shah I_d vs V_ds
.include CMOS.txt


v_dd 1 0 3.3
v_in 2 0 pulse(0 3.3 0 20p 20p 280p 600p)
v_bb_p 10 0 3.3
v_bb_n 11 0 0

m_p 3 2 1 10 cmosp L=0.4u W=3.36u
m_n 3 2 0 11 cmosn L=0.4u W=1.3u
c0 3 4 0.05p
v_dummy 4 0 0

.tran 0.1p 5000p
.control
run
meas tran rise trig v(3) val=0.33 rise=1 targ v(3) val=2.97 rise=1
meas tran delay trig v(2) val=1.665 rise=2 targ v(3) val=1.665 fall=2
meas tran fall trig v(3) val=2.97 fall=1 targ v(3) val=0.33 fall=1

.endc
.end