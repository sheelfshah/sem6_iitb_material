19D070052 Sheel Shah Solar IV
.include Solar_Cell.txt

r2 0 22 100
x2 22 32 solar_cell IL_val = 8e-3
v_dummy2 0 32 0

r3 0 23 100
x3 23 33 solar_cell IL_val = 10e-3
v_dummy3 0 33 0
** 1: dark, 2: 8mA, 3: 10mA
* start control
.control
set color0 = rgb:f/f/e
set color1 = rgb:1/1/1

run

dc r2 1 500 1
let i1 = i(v_dummy2)
let v1 = v(22)-v(32)
let p1 = i1*v1

dc r3 1 500 1
plot dc1.i1 vs dc1.v1, i(v_dummy3) vs v(23)-v(33)
plot dc1.p1 vs dc1.v1, i(v_dummy3)*(v(23)-v(33)) vs v(23)-v(33)

** i_sc1 = 7.9mA, i_sc2 = 9.9mA
** v_oc1 = 411.6mV, v_oc2 = 425.3mV
** v_mp1 = 278mV, p_mp1 = 1.73mW
** v_mp2 = 278.6mV, p_mp2 = 2.15mW
** ff1 = 0.53
** ff2 = 0.51
* end control
.endc

.end