19D070052 Sheel Shah I_d vs V_ds

.include NMOSFET.txt

** 1 2 3 4: drain gate source body
m_short 11 2 0 4 NMOSFET W=1.2u L=0.2u
m_long 12 2 0 4 NMOSFET W=120u L=20u
v_dd 4 0 0
v_id1 10 11 0
v_id2 10 12 0
v_ds 10 0 3
v_gs 2 0


.dc v_gs 0 3.3 0.01

* start control
.control
run
 
plot i(v_id1), i(v_id2) vs v(2)
plot log10(i(v_id1)), log10(i(v_id2)) vs v(2)

** v_th: 0.1V, 0.5V
** i_on: 1.47m, 2.45m
** ss: 166mV/dec, 104mV/dec
** i_off: 2e-6, 6.3e-12

** ro: 41k, 1300k

.endc

.end