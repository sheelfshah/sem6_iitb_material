Sheel Shah 19D070052

.include bc547.txt

q0 2 0 1 bc547a
r1 1 3 100
v2 3 0
i_e 2 0

.dc v2  -3.5 100 0.1 i_e 0 10m 1m

.control
run
plot  -i(v2) vs v(1)

.endc
.end
