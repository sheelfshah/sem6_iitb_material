19d070052 rf switch

.include rn142s.txt
.include Diode_1N914.txt

v_in 1 0 sin(0 3 10000k 0 0)
c1 1 2 100n
r1 2 0 500
v_diode 2 21 0
d_diode 21 3 1N914
r2 3 4 500
v_bias 4 0 5
c2 3 51 100n
v_out 51 5 0
r3 5 0 50

.tran 1n 0.5u
.control

run
plot v(5) v(1)
.endc

.end