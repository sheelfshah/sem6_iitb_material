Sheel Shah 19D070052

.include bc547a.txt

q0 0 1 2 bc547a
r2 3 2 100
i_source 0 1 0.1m
v_ce 3 0 pulse(0 3 0 0 0 0.25u 1000)

.tran 1n 1u
.control
run

plot -i(v_ce)
** time = 1e-8

.endc
.end 
