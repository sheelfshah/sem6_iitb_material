19D070052 Sheel Shah IV

.include Diode_1N914.txt
.include BZT52C18S.txt

v_dc 1 0

* r11 1 21 100
* r21 21 0 1k
* v_d1 21 31 0
* d01 31 41 1N914
* r31 41 0 100

r12 1 22 100
r22 22 0 1k
v_d2 22 32 0
x02 42 32 DI_BZT52C18S
r32 42 0 100

.dc v_dc -3 0 0.01 temp 20 30 10

.control

run

* plot i(v_d1) vs v(31)-v(41), (2m) vs v(31)-v(41)
plot i(v_d2) vs v(32)-v(42), (-0.5m) vs v(32)-v(42)

.endc

.end

** v_d pn: (20 to 80), i = 2m
** 0.655, 0.637, 0.618, 0.600, 0.582, 0.563, 0.544
** slope = -1.85 mV/C

** v_d zen: (20 to 80), i = -0.5m
** -0.556, -0.534, -0.512, -0.490, -0.468, -0.445, -0.422
** slope = 2.23 mV/C