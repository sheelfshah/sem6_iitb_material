19D070052 Sheel Shah I_d vs V_ds
.include PMOS_NMOS.txt


v_dd 1 0 3.3
v_in 2 0 pulse(0 3.3v 0 500p 500p 4500p 10n)
v_bb_p 10 0 3
v_bb_n 11 0 0.3

m_p 3 2 1 10 cmosp L=0.4u W=2.9u AS=4.8e-11 PS=121.6u AD=4.8e-11 PD=121.6u
m_n 3 2 0 11 cmosn L=0.4u W=1.2u
c0 3 4 200f
v_dummy 4 0 0

.tran 2p 40n
.control
run
meas tran rise trig v(3) val=0.33 rise=1 targ v(3) val=2.97 rise=1
meas tran delay trig v(2) val=1.665 rise=2 targ v(3) val=1.665 fall=2
meas tran fall trig v(3) val=2.97 fall=1 targ v(3) val=0.33 fall=1
meas tran i_peak_charging MAX i(v_dummy)
meas tran i_peak_charging MIN i(v_dummy)


** table
** bb_n, bb_p, pcc, pdc, dt
** 0.3, 3, 6.07e-4, -4.76e-4, 7.94e-10
** 0.1, 3.2, 6.07e-4, -4.80e-4m, 7.88e-10
** 0, 3.3, 6.04e-4, -4.79e-4, 7.89e-10
** -0.5, 3.8, 5.87e-4, -4.74e-4, 8.00e-10
** -1, 4.3, 5.72e-4, -4.71 e-4, 8.11e-10


** as v_b changes, v_t changes, and hence i_ds changes.
** as bb_p increases, thresh_p increases, i_ds_p decreases (curve shifts to left)
** similarly i_ds_n decreases in magnitude too

** delay is higher when body bias is applied
** v_th_n/v_th_p decreases as bb is increased and vice versa

** case 5 as it has lowest capacitor currents
.endc
.end